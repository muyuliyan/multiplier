//unsigned num multipiler

module mult_gen_1(
    input CLK,
    input mul,
    input [31:0] A,
    input [31:0] B,
    output [63:0] P,
    input SCLR,
);
