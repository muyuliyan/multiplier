/*a 2 bit booth wallace tree multiplier*/

module multipiler(
    input mul_clk,
    input resetn,
    input mul_signed,
    input [31:0]x,
    input [31:0]y,
    output [63:0]result
);






endmodule


.Inu1-C1k（mu1-C1k）′
.rese仁n（resetn）′
ˉmu1-s1gned（mu1-signed）′
。×（×）〃
.y（y）′
.reSu1仁（reSu1t）
