//signed num multiplier

module mult_gen_0(
    input CLK,
    input [31:0]A,
    input [31:0]B,
    output [31:0]P,
    input SCLR,
)
